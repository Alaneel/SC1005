module main(input A, B, X, Y, output Out);

    assign Out = (A > B) ? X : Y;

endmodule